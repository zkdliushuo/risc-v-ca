
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h8492acf5;
    ram_cell[       1] = 32'h0;  // 32'h9d0f8dcc;
    ram_cell[       2] = 32'h0;  // 32'hbd889cda;
    ram_cell[       3] = 32'h0;  // 32'h3266cbb4;
    ram_cell[       4] = 32'h0;  // 32'hbe28e36a;
    ram_cell[       5] = 32'h0;  // 32'h7591f2f7;
    ram_cell[       6] = 32'h0;  // 32'h3fc3b6fa;
    ram_cell[       7] = 32'h0;  // 32'hb709d4b7;
    ram_cell[       8] = 32'h0;  // 32'hed3b8f96;
    ram_cell[       9] = 32'h0;  // 32'h3dc1bca3;
    ram_cell[      10] = 32'h0;  // 32'h5499e9cd;
    ram_cell[      11] = 32'h0;  // 32'hf7804622;
    ram_cell[      12] = 32'h0;  // 32'hff1438c7;
    ram_cell[      13] = 32'h0;  // 32'h7b1e7dc1;
    ram_cell[      14] = 32'h0;  // 32'h0beea247;
    ram_cell[      15] = 32'h0;  // 32'h7f511a8e;
    ram_cell[      16] = 32'h0;  // 32'he610643e;
    ram_cell[      17] = 32'h0;  // 32'h5747e9f4;
    ram_cell[      18] = 32'h0;  // 32'h6c8bfc0a;
    ram_cell[      19] = 32'h0;  // 32'hd537de26;
    ram_cell[      20] = 32'h0;  // 32'h08dfe84d;
    ram_cell[      21] = 32'h0;  // 32'h1fd10544;
    ram_cell[      22] = 32'h0;  // 32'h9f5693d4;
    ram_cell[      23] = 32'h0;  // 32'hb1950c83;
    ram_cell[      24] = 32'h0;  // 32'h5f2afca1;
    ram_cell[      25] = 32'h0;  // 32'h8ed201d3;
    ram_cell[      26] = 32'h0;  // 32'h11b8790f;
    ram_cell[      27] = 32'h0;  // 32'h4762249a;
    ram_cell[      28] = 32'h0;  // 32'hee547816;
    ram_cell[      29] = 32'h0;  // 32'h8f11e516;
    ram_cell[      30] = 32'h0;  // 32'he3fb08aa;
    ram_cell[      31] = 32'h0;  // 32'h8d5c409e;
    ram_cell[      32] = 32'h0;  // 32'hcf88a103;
    ram_cell[      33] = 32'h0;  // 32'h151de1d2;
    ram_cell[      34] = 32'h0;  // 32'hb9544e63;
    ram_cell[      35] = 32'h0;  // 32'hbd762a95;
    ram_cell[      36] = 32'h0;  // 32'h019becd5;
    ram_cell[      37] = 32'h0;  // 32'h87bdb738;
    ram_cell[      38] = 32'h0;  // 32'h4ebc2ec0;
    ram_cell[      39] = 32'h0;  // 32'hf39741d3;
    ram_cell[      40] = 32'h0;  // 32'h4782cd30;
    ram_cell[      41] = 32'h0;  // 32'he2cce973;
    ram_cell[      42] = 32'h0;  // 32'hed6ae67d;
    ram_cell[      43] = 32'h0;  // 32'h8cd15b3e;
    ram_cell[      44] = 32'h0;  // 32'ha64d828f;
    ram_cell[      45] = 32'h0;  // 32'h1ba8f315;
    ram_cell[      46] = 32'h0;  // 32'h26dab35e;
    ram_cell[      47] = 32'h0;  // 32'h868c54b2;
    ram_cell[      48] = 32'h0;  // 32'heaacddae;
    ram_cell[      49] = 32'h0;  // 32'h9dcfba7b;
    ram_cell[      50] = 32'h0;  // 32'head2e7c7;
    ram_cell[      51] = 32'h0;  // 32'h6df0b15a;
    ram_cell[      52] = 32'h0;  // 32'h2eced7ee;
    ram_cell[      53] = 32'h0;  // 32'h19f9a627;
    ram_cell[      54] = 32'h0;  // 32'h02b36a6f;
    ram_cell[      55] = 32'h0;  // 32'h02285299;
    ram_cell[      56] = 32'h0;  // 32'h81d0cdee;
    ram_cell[      57] = 32'h0;  // 32'h1339efff;
    ram_cell[      58] = 32'h0;  // 32'ha82629d6;
    ram_cell[      59] = 32'h0;  // 32'ha1668e01;
    ram_cell[      60] = 32'h0;  // 32'h8b882051;
    ram_cell[      61] = 32'h0;  // 32'h5d4ac4d5;
    ram_cell[      62] = 32'h0;  // 32'h06254cd5;
    ram_cell[      63] = 32'h0;  // 32'h2ccf3d1e;
    ram_cell[      64] = 32'h0;  // 32'h6f37c989;
    ram_cell[      65] = 32'h0;  // 32'h8bc2ddaf;
    ram_cell[      66] = 32'h0;  // 32'hcd16b02c;
    ram_cell[      67] = 32'h0;  // 32'h267d67b7;
    ram_cell[      68] = 32'h0;  // 32'h7a90ac4d;
    ram_cell[      69] = 32'h0;  // 32'h9f3e0277;
    ram_cell[      70] = 32'h0;  // 32'hc0ccd788;
    ram_cell[      71] = 32'h0;  // 32'h6746b7d2;
    ram_cell[      72] = 32'h0;  // 32'h51cc888a;
    ram_cell[      73] = 32'h0;  // 32'haafe0d5c;
    ram_cell[      74] = 32'h0;  // 32'h70eeabcd;
    ram_cell[      75] = 32'h0;  // 32'h0cc10bf2;
    ram_cell[      76] = 32'h0;  // 32'h8a0b3df8;
    ram_cell[      77] = 32'h0;  // 32'hc3489792;
    ram_cell[      78] = 32'h0;  // 32'hf9bb70ca;
    ram_cell[      79] = 32'h0;  // 32'hb9587d69;
    ram_cell[      80] = 32'h0;  // 32'h2c6b6386;
    ram_cell[      81] = 32'h0;  // 32'h4590c01b;
    ram_cell[      82] = 32'h0;  // 32'h9888ec9c;
    ram_cell[      83] = 32'h0;  // 32'h71a61038;
    ram_cell[      84] = 32'h0;  // 32'h80eb9772;
    ram_cell[      85] = 32'h0;  // 32'h13a3bac3;
    ram_cell[      86] = 32'h0;  // 32'h661da566;
    ram_cell[      87] = 32'h0;  // 32'he4fb028f;
    ram_cell[      88] = 32'h0;  // 32'h87787ddb;
    ram_cell[      89] = 32'h0;  // 32'h5e026014;
    ram_cell[      90] = 32'h0;  // 32'hf399a392;
    ram_cell[      91] = 32'h0;  // 32'h8a763a5b;
    ram_cell[      92] = 32'h0;  // 32'h8e667253;
    ram_cell[      93] = 32'h0;  // 32'hcedd5c22;
    ram_cell[      94] = 32'h0;  // 32'hf871edee;
    ram_cell[      95] = 32'h0;  // 32'h000b5b15;
    ram_cell[      96] = 32'h0;  // 32'h7c3aa757;
    ram_cell[      97] = 32'h0;  // 32'h9468cc6b;
    ram_cell[      98] = 32'h0;  // 32'hfcad75f2;
    ram_cell[      99] = 32'h0;  // 32'hb1f1f0f7;
    ram_cell[     100] = 32'h0;  // 32'h7ecfb0ed;
    ram_cell[     101] = 32'h0;  // 32'h06830a79;
    ram_cell[     102] = 32'h0;  // 32'hce68f1a1;
    ram_cell[     103] = 32'h0;  // 32'hd7dd5e5c;
    ram_cell[     104] = 32'h0;  // 32'h853270e3;
    ram_cell[     105] = 32'h0;  // 32'hc873fdc4;
    ram_cell[     106] = 32'h0;  // 32'hf417bdbc;
    ram_cell[     107] = 32'h0;  // 32'h6dd6d049;
    ram_cell[     108] = 32'h0;  // 32'h0e33adc7;
    ram_cell[     109] = 32'h0;  // 32'hba85d720;
    ram_cell[     110] = 32'h0;  // 32'h032d3ba8;
    ram_cell[     111] = 32'h0;  // 32'h6ee45515;
    ram_cell[     112] = 32'h0;  // 32'h4d36fa21;
    ram_cell[     113] = 32'h0;  // 32'h8b39d59e;
    ram_cell[     114] = 32'h0;  // 32'h8982d6de;
    ram_cell[     115] = 32'h0;  // 32'hfa172b82;
    ram_cell[     116] = 32'h0;  // 32'h702b4603;
    ram_cell[     117] = 32'h0;  // 32'he58afbc7;
    ram_cell[     118] = 32'h0;  // 32'hdb9bb0df;
    ram_cell[     119] = 32'h0;  // 32'h4760ed1b;
    ram_cell[     120] = 32'h0;  // 32'h1681e3c3;
    ram_cell[     121] = 32'h0;  // 32'h4edfec9c;
    ram_cell[     122] = 32'h0;  // 32'hd0c09e78;
    ram_cell[     123] = 32'h0;  // 32'h19158844;
    ram_cell[     124] = 32'h0;  // 32'hdacfae4c;
    ram_cell[     125] = 32'h0;  // 32'hde10047e;
    ram_cell[     126] = 32'h0;  // 32'heb79c2e8;
    ram_cell[     127] = 32'h0;  // 32'h599a7e45;
    ram_cell[     128] = 32'h0;  // 32'h1ad0c5f4;
    ram_cell[     129] = 32'h0;  // 32'hf83073b6;
    ram_cell[     130] = 32'h0;  // 32'h45a71179;
    ram_cell[     131] = 32'h0;  // 32'h2587fc7d;
    ram_cell[     132] = 32'h0;  // 32'hccf561d9;
    ram_cell[     133] = 32'h0;  // 32'h98a82a32;
    ram_cell[     134] = 32'h0;  // 32'h56c42e85;
    ram_cell[     135] = 32'h0;  // 32'h0fb6bfb1;
    ram_cell[     136] = 32'h0;  // 32'h97ee156d;
    ram_cell[     137] = 32'h0;  // 32'h6320eae1;
    ram_cell[     138] = 32'h0;  // 32'hcbc0e8b9;
    ram_cell[     139] = 32'h0;  // 32'h9dc9c165;
    ram_cell[     140] = 32'h0;  // 32'hee7eea59;
    ram_cell[     141] = 32'h0;  // 32'h1d1335d6;
    ram_cell[     142] = 32'h0;  // 32'hfd83d785;
    ram_cell[     143] = 32'h0;  // 32'h60eb6cab;
    ram_cell[     144] = 32'h0;  // 32'hbdc4474d;
    ram_cell[     145] = 32'h0;  // 32'hcaa6f6b0;
    ram_cell[     146] = 32'h0;  // 32'hdceacfe9;
    ram_cell[     147] = 32'h0;  // 32'h5a1c5354;
    ram_cell[     148] = 32'h0;  // 32'h9646d0d8;
    ram_cell[     149] = 32'h0;  // 32'h5ea7dbc1;
    ram_cell[     150] = 32'h0;  // 32'hb96b1e7c;
    ram_cell[     151] = 32'h0;  // 32'h02d4f324;
    ram_cell[     152] = 32'h0;  // 32'h43728b4f;
    ram_cell[     153] = 32'h0;  // 32'h3939088c;
    ram_cell[     154] = 32'h0;  // 32'h25a576dc;
    ram_cell[     155] = 32'h0;  // 32'h4cc507f4;
    ram_cell[     156] = 32'h0;  // 32'hc227f0fa;
    ram_cell[     157] = 32'h0;  // 32'h3839e30f;
    ram_cell[     158] = 32'h0;  // 32'h2081c962;
    ram_cell[     159] = 32'h0;  // 32'hcd0cf4e8;
    ram_cell[     160] = 32'h0;  // 32'h9b1b1432;
    ram_cell[     161] = 32'h0;  // 32'h2d6f6a68;
    ram_cell[     162] = 32'h0;  // 32'h88862fb3;
    ram_cell[     163] = 32'h0;  // 32'h44389a2d;
    ram_cell[     164] = 32'h0;  // 32'hcc02faca;
    ram_cell[     165] = 32'h0;  // 32'h5ea8df0e;
    ram_cell[     166] = 32'h0;  // 32'h40a81690;
    ram_cell[     167] = 32'h0;  // 32'h5eefcb32;
    ram_cell[     168] = 32'h0;  // 32'h589aba63;
    ram_cell[     169] = 32'h0;  // 32'hf6b6fb1d;
    ram_cell[     170] = 32'h0;  // 32'hc3ae66d9;
    ram_cell[     171] = 32'h0;  // 32'hb0f312a8;
    ram_cell[     172] = 32'h0;  // 32'hedfa6844;
    ram_cell[     173] = 32'h0;  // 32'hd0dbe00e;
    ram_cell[     174] = 32'h0;  // 32'heb3809c9;
    ram_cell[     175] = 32'h0;  // 32'h9986bfa0;
    ram_cell[     176] = 32'h0;  // 32'h6af05d94;
    ram_cell[     177] = 32'h0;  // 32'ha3f7f106;
    ram_cell[     178] = 32'h0;  // 32'h0627fcb9;
    ram_cell[     179] = 32'h0;  // 32'h9e569af8;
    ram_cell[     180] = 32'h0;  // 32'hb4872ff4;
    ram_cell[     181] = 32'h0;  // 32'hee94c63d;
    ram_cell[     182] = 32'h0;  // 32'hd97399aa;
    ram_cell[     183] = 32'h0;  // 32'he075deb2;
    ram_cell[     184] = 32'h0;  // 32'he65f2054;
    ram_cell[     185] = 32'h0;  // 32'ha80df28e;
    ram_cell[     186] = 32'h0;  // 32'ha729307f;
    ram_cell[     187] = 32'h0;  // 32'h65846871;
    ram_cell[     188] = 32'h0;  // 32'h68dccfd7;
    ram_cell[     189] = 32'h0;  // 32'hc458eb67;
    ram_cell[     190] = 32'h0;  // 32'h372844c9;
    ram_cell[     191] = 32'h0;  // 32'h3b3f8ce8;
    ram_cell[     192] = 32'h0;  // 32'h9bb35f90;
    ram_cell[     193] = 32'h0;  // 32'h98ba11f4;
    ram_cell[     194] = 32'h0;  // 32'h11135bc0;
    ram_cell[     195] = 32'h0;  // 32'h443298ca;
    ram_cell[     196] = 32'h0;  // 32'hb048318f;
    ram_cell[     197] = 32'h0;  // 32'h6ee1f3c0;
    ram_cell[     198] = 32'h0;  // 32'h2196eda3;
    ram_cell[     199] = 32'h0;  // 32'h535bcf82;
    ram_cell[     200] = 32'h0;  // 32'h36c965bf;
    ram_cell[     201] = 32'h0;  // 32'he285f898;
    ram_cell[     202] = 32'h0;  // 32'he4422091;
    ram_cell[     203] = 32'h0;  // 32'hb2ec33ee;
    ram_cell[     204] = 32'h0;  // 32'hbae62c5c;
    ram_cell[     205] = 32'h0;  // 32'hf74a433d;
    ram_cell[     206] = 32'h0;  // 32'ha9034809;
    ram_cell[     207] = 32'h0;  // 32'hfbed9c27;
    ram_cell[     208] = 32'h0;  // 32'h572316f9;
    ram_cell[     209] = 32'h0;  // 32'h56bb56ca;
    ram_cell[     210] = 32'h0;  // 32'h5c73fa29;
    ram_cell[     211] = 32'h0;  // 32'h46a57f8b;
    ram_cell[     212] = 32'h0;  // 32'h0ddad7ad;
    ram_cell[     213] = 32'h0;  // 32'h5614850e;
    ram_cell[     214] = 32'h0;  // 32'h1d9bb52d;
    ram_cell[     215] = 32'h0;  // 32'hc232fcfb;
    ram_cell[     216] = 32'h0;  // 32'ha69cefd2;
    ram_cell[     217] = 32'h0;  // 32'h994092ba;
    ram_cell[     218] = 32'h0;  // 32'h5ebb31e4;
    ram_cell[     219] = 32'h0;  // 32'h18fa9d87;
    ram_cell[     220] = 32'h0;  // 32'h80852829;
    ram_cell[     221] = 32'h0;  // 32'hb08aef95;
    ram_cell[     222] = 32'h0;  // 32'h50b98a44;
    ram_cell[     223] = 32'h0;  // 32'h4537e19f;
    ram_cell[     224] = 32'h0;  // 32'hdb001110;
    ram_cell[     225] = 32'h0;  // 32'hd9f23349;
    ram_cell[     226] = 32'h0;  // 32'h17d4785e;
    ram_cell[     227] = 32'h0;  // 32'h717e94af;
    ram_cell[     228] = 32'h0;  // 32'h009d49a5;
    ram_cell[     229] = 32'h0;  // 32'h1dd75ab6;
    ram_cell[     230] = 32'h0;  // 32'h908cc6c8;
    ram_cell[     231] = 32'h0;  // 32'h3a8cfc77;
    ram_cell[     232] = 32'h0;  // 32'he87bb95a;
    ram_cell[     233] = 32'h0;  // 32'hcf2bd61e;
    ram_cell[     234] = 32'h0;  // 32'h315979c9;
    ram_cell[     235] = 32'h0;  // 32'h1b56bd08;
    ram_cell[     236] = 32'h0;  // 32'h2bd63696;
    ram_cell[     237] = 32'h0;  // 32'hd8701944;
    ram_cell[     238] = 32'h0;  // 32'h08c13fc4;
    ram_cell[     239] = 32'h0;  // 32'hc85db988;
    ram_cell[     240] = 32'h0;  // 32'h2f3c49e0;
    ram_cell[     241] = 32'h0;  // 32'h3a23144d;
    ram_cell[     242] = 32'h0;  // 32'h62816a0c;
    ram_cell[     243] = 32'h0;  // 32'h07dd9de9;
    ram_cell[     244] = 32'h0;  // 32'hf83f843b;
    ram_cell[     245] = 32'h0;  // 32'hf0ecdfd9;
    ram_cell[     246] = 32'h0;  // 32'hf2a95d52;
    ram_cell[     247] = 32'h0;  // 32'h79655b26;
    ram_cell[     248] = 32'h0;  // 32'hfe69d7a8;
    ram_cell[     249] = 32'h0;  // 32'hd6a8d1a1;
    ram_cell[     250] = 32'h0;  // 32'hf8b76553;
    ram_cell[     251] = 32'h0;  // 32'h3ce91869;
    ram_cell[     252] = 32'h0;  // 32'h7cacdb93;
    ram_cell[     253] = 32'h0;  // 32'hc9d7149a;
    ram_cell[     254] = 32'h0;  // 32'hf751c75c;
    ram_cell[     255] = 32'h0;  // 32'h78e341e6;
    // src matrix A
    ram_cell[     256] = 32'h9638b9e1;
    ram_cell[     257] = 32'ha36e633b;
    ram_cell[     258] = 32'h21514ec1;
    ram_cell[     259] = 32'hdca3a564;
    ram_cell[     260] = 32'h9703112e;
    ram_cell[     261] = 32'heed843e0;
    ram_cell[     262] = 32'h8a77a92c;
    ram_cell[     263] = 32'hd72cbc30;
    ram_cell[     264] = 32'he79b369a;
    ram_cell[     265] = 32'h28b79c10;
    ram_cell[     266] = 32'h76285265;
    ram_cell[     267] = 32'hd54a3fc6;
    ram_cell[     268] = 32'h9c8caff9;
    ram_cell[     269] = 32'hfad60df4;
    ram_cell[     270] = 32'hded4058f;
    ram_cell[     271] = 32'h82ad726e;
    ram_cell[     272] = 32'h444b0653;
    ram_cell[     273] = 32'h0ea3ae4a;
    ram_cell[     274] = 32'h81bec1af;
    ram_cell[     275] = 32'hf8c79ea9;
    ram_cell[     276] = 32'h98ab56a2;
    ram_cell[     277] = 32'hb6db8df9;
    ram_cell[     278] = 32'he19fc651;
    ram_cell[     279] = 32'h3d67401b;
    ram_cell[     280] = 32'h137c95b0;
    ram_cell[     281] = 32'h4ebbeda2;
    ram_cell[     282] = 32'h3a72e1e2;
    ram_cell[     283] = 32'ha2193600;
    ram_cell[     284] = 32'hbc09ed72;
    ram_cell[     285] = 32'hf1140a0c;
    ram_cell[     286] = 32'h1b4d29d6;
    ram_cell[     287] = 32'h13d080c5;
    ram_cell[     288] = 32'h282f2eb0;
    ram_cell[     289] = 32'h025cbaa0;
    ram_cell[     290] = 32'h14cfea8d;
    ram_cell[     291] = 32'h048e45d0;
    ram_cell[     292] = 32'h6a6d3409;
    ram_cell[     293] = 32'h819b737e;
    ram_cell[     294] = 32'h617d240a;
    ram_cell[     295] = 32'h91093110;
    ram_cell[     296] = 32'h77361350;
    ram_cell[     297] = 32'h0937aeef;
    ram_cell[     298] = 32'h6a06f745;
    ram_cell[     299] = 32'h9a0ebd1f;
    ram_cell[     300] = 32'h84ff5238;
    ram_cell[     301] = 32'hba5db3b3;
    ram_cell[     302] = 32'hea093aef;
    ram_cell[     303] = 32'hb8a2c635;
    ram_cell[     304] = 32'h62377279;
    ram_cell[     305] = 32'h96cb8322;
    ram_cell[     306] = 32'h4eb36d0a;
    ram_cell[     307] = 32'h63b02fa4;
    ram_cell[     308] = 32'h72a52db6;
    ram_cell[     309] = 32'h2aa6371c;
    ram_cell[     310] = 32'h88206d7a;
    ram_cell[     311] = 32'h48210787;
    ram_cell[     312] = 32'ha6daf7f6;
    ram_cell[     313] = 32'h23a59365;
    ram_cell[     314] = 32'h05d6bd52;
    ram_cell[     315] = 32'ha6c38158;
    ram_cell[     316] = 32'h365542cc;
    ram_cell[     317] = 32'h2c6f73de;
    ram_cell[     318] = 32'hfb02059c;
    ram_cell[     319] = 32'h36aef1cb;
    ram_cell[     320] = 32'hec713b0d;
    ram_cell[     321] = 32'hf216ce16;
    ram_cell[     322] = 32'heaa5dafd;
    ram_cell[     323] = 32'h682f4726;
    ram_cell[     324] = 32'h746316a7;
    ram_cell[     325] = 32'h467fed5a;
    ram_cell[     326] = 32'he4f9ffa3;
    ram_cell[     327] = 32'hc47305b5;
    ram_cell[     328] = 32'hf3339336;
    ram_cell[     329] = 32'h63bfa4f4;
    ram_cell[     330] = 32'hc7deeb94;
    ram_cell[     331] = 32'h6fda254c;
    ram_cell[     332] = 32'he32774ca;
    ram_cell[     333] = 32'h08a6211a;
    ram_cell[     334] = 32'h957af49d;
    ram_cell[     335] = 32'h9a088a1a;
    ram_cell[     336] = 32'hdbba299c;
    ram_cell[     337] = 32'h59bf2486;
    ram_cell[     338] = 32'he1309f08;
    ram_cell[     339] = 32'h6219013c;
    ram_cell[     340] = 32'hece8ee4a;
    ram_cell[     341] = 32'h394a6f3a;
    ram_cell[     342] = 32'hf4aa32c4;
    ram_cell[     343] = 32'h580df057;
    ram_cell[     344] = 32'h032256c9;
    ram_cell[     345] = 32'h5c0efff8;
    ram_cell[     346] = 32'h1eac31cc;
    ram_cell[     347] = 32'h95b70e08;
    ram_cell[     348] = 32'hba5a822e;
    ram_cell[     349] = 32'hc1b9802f;
    ram_cell[     350] = 32'h4de4e0a0;
    ram_cell[     351] = 32'h13361819;
    ram_cell[     352] = 32'h7e713955;
    ram_cell[     353] = 32'h437938c3;
    ram_cell[     354] = 32'h1598601c;
    ram_cell[     355] = 32'h70823ee7;
    ram_cell[     356] = 32'h34d9593a;
    ram_cell[     357] = 32'h2e850b54;
    ram_cell[     358] = 32'h46420ec8;
    ram_cell[     359] = 32'h1d15b75a;
    ram_cell[     360] = 32'h70893486;
    ram_cell[     361] = 32'h03f1640e;
    ram_cell[     362] = 32'hdf7fdae8;
    ram_cell[     363] = 32'ha5e3ebe5;
    ram_cell[     364] = 32'hdbc653bf;
    ram_cell[     365] = 32'h4189958a;
    ram_cell[     366] = 32'hbe1e87f5;
    ram_cell[     367] = 32'hfc5ff20b;
    ram_cell[     368] = 32'h2b24c427;
    ram_cell[     369] = 32'haa798ef8;
    ram_cell[     370] = 32'h1b7f199a;
    ram_cell[     371] = 32'ha1af65ce;
    ram_cell[     372] = 32'hd497c186;
    ram_cell[     373] = 32'h926688fd;
    ram_cell[     374] = 32'hc4422f07;
    ram_cell[     375] = 32'hbac39ee6;
    ram_cell[     376] = 32'hfc16d172;
    ram_cell[     377] = 32'h102fdb8b;
    ram_cell[     378] = 32'h64edae94;
    ram_cell[     379] = 32'h1cdee50f;
    ram_cell[     380] = 32'h2f7fd178;
    ram_cell[     381] = 32'h028fbd53;
    ram_cell[     382] = 32'h15706f2a;
    ram_cell[     383] = 32'h5004a39d;
    ram_cell[     384] = 32'h0ff9f131;
    ram_cell[     385] = 32'hefd30340;
    ram_cell[     386] = 32'hedd5c5cb;
    ram_cell[     387] = 32'h517e8c9f;
    ram_cell[     388] = 32'h998984ae;
    ram_cell[     389] = 32'h9a4a2a63;
    ram_cell[     390] = 32'hb537de39;
    ram_cell[     391] = 32'h552c4c0e;
    ram_cell[     392] = 32'hff08d7b2;
    ram_cell[     393] = 32'h8f280dfd;
    ram_cell[     394] = 32'h13b474ef;
    ram_cell[     395] = 32'h5005626f;
    ram_cell[     396] = 32'hafd80fc3;
    ram_cell[     397] = 32'h9fe4549d;
    ram_cell[     398] = 32'hc075f395;
    ram_cell[     399] = 32'h6b391321;
    ram_cell[     400] = 32'h9ea3f628;
    ram_cell[     401] = 32'hb329032b;
    ram_cell[     402] = 32'h71c8fba4;
    ram_cell[     403] = 32'h73b2b2f9;
    ram_cell[     404] = 32'h49de4475;
    ram_cell[     405] = 32'h33b22095;
    ram_cell[     406] = 32'h9610ab14;
    ram_cell[     407] = 32'h41c02e0f;
    ram_cell[     408] = 32'h0b101006;
    ram_cell[     409] = 32'hc0e4155d;
    ram_cell[     410] = 32'hc88a9862;
    ram_cell[     411] = 32'h4aa409c6;
    ram_cell[     412] = 32'hb64cd5bc;
    ram_cell[     413] = 32'hb2bfc594;
    ram_cell[     414] = 32'h990a4324;
    ram_cell[     415] = 32'hcadcbb30;
    ram_cell[     416] = 32'h4379a99d;
    ram_cell[     417] = 32'h9e2a5701;
    ram_cell[     418] = 32'h1a65d9d1;
    ram_cell[     419] = 32'h5e838483;
    ram_cell[     420] = 32'hb7a7fb27;
    ram_cell[     421] = 32'ha10268fb;
    ram_cell[     422] = 32'hab731b5e;
    ram_cell[     423] = 32'hfc07d697;
    ram_cell[     424] = 32'he9596bdb;
    ram_cell[     425] = 32'he0aa0a60;
    ram_cell[     426] = 32'h75ad1e2e;
    ram_cell[     427] = 32'h893601b6;
    ram_cell[     428] = 32'h659956d0;
    ram_cell[     429] = 32'hcac64961;
    ram_cell[     430] = 32'h6e9ae393;
    ram_cell[     431] = 32'hb9166f70;
    ram_cell[     432] = 32'h08060938;
    ram_cell[     433] = 32'h742afc71;
    ram_cell[     434] = 32'hd99b75b1;
    ram_cell[     435] = 32'h936eea7d;
    ram_cell[     436] = 32'h50824a76;
    ram_cell[     437] = 32'hd99ebb75;
    ram_cell[     438] = 32'h63b8a65d;
    ram_cell[     439] = 32'h7af41812;
    ram_cell[     440] = 32'hd352347e;
    ram_cell[     441] = 32'h30943c02;
    ram_cell[     442] = 32'h1390162e;
    ram_cell[     443] = 32'h3dc0a9f1;
    ram_cell[     444] = 32'h2170533a;
    ram_cell[     445] = 32'h4559ac0f;
    ram_cell[     446] = 32'hc4a6efe5;
    ram_cell[     447] = 32'h92ec4201;
    ram_cell[     448] = 32'h429baa38;
    ram_cell[     449] = 32'hb8da6b10;
    ram_cell[     450] = 32'h78557747;
    ram_cell[     451] = 32'hfa3d5519;
    ram_cell[     452] = 32'h7a10bd19;
    ram_cell[     453] = 32'h26a0ca01;
    ram_cell[     454] = 32'h75b82d10;
    ram_cell[     455] = 32'h407c2237;
    ram_cell[     456] = 32'hcfd139b8;
    ram_cell[     457] = 32'h2cfcdab1;
    ram_cell[     458] = 32'h8ebceaa4;
    ram_cell[     459] = 32'hb830feb8;
    ram_cell[     460] = 32'hc33ad727;
    ram_cell[     461] = 32'h7d2986c4;
    ram_cell[     462] = 32'haab037de;
    ram_cell[     463] = 32'hae2f3415;
    ram_cell[     464] = 32'h4dc7bbe1;
    ram_cell[     465] = 32'hd76d2413;
    ram_cell[     466] = 32'ha602dc71;
    ram_cell[     467] = 32'hb68c9b69;
    ram_cell[     468] = 32'h32a45789;
    ram_cell[     469] = 32'he1f9b3a2;
    ram_cell[     470] = 32'h1dde00e7;
    ram_cell[     471] = 32'h2d463f3d;
    ram_cell[     472] = 32'hb32574d6;
    ram_cell[     473] = 32'hb3959a08;
    ram_cell[     474] = 32'hb1aafe73;
    ram_cell[     475] = 32'he47925cf;
    ram_cell[     476] = 32'h40fccdac;
    ram_cell[     477] = 32'h51d93831;
    ram_cell[     478] = 32'h2bbff1b6;
    ram_cell[     479] = 32'hdb23b9d3;
    ram_cell[     480] = 32'h02744627;
    ram_cell[     481] = 32'h8932190e;
    ram_cell[     482] = 32'h14f129bc;
    ram_cell[     483] = 32'h6b907dc4;
    ram_cell[     484] = 32'h93fb1a6f;
    ram_cell[     485] = 32'had004461;
    ram_cell[     486] = 32'h4908de53;
    ram_cell[     487] = 32'h76dbe5d0;
    ram_cell[     488] = 32'h1d416f52;
    ram_cell[     489] = 32'hebff8371;
    ram_cell[     490] = 32'h286e3016;
    ram_cell[     491] = 32'h7d5b889d;
    ram_cell[     492] = 32'h3cb2afa9;
    ram_cell[     493] = 32'heb8197a0;
    ram_cell[     494] = 32'h5432ef09;
    ram_cell[     495] = 32'hc2c3982d;
    ram_cell[     496] = 32'h1d2df6c1;
    ram_cell[     497] = 32'h572e48ac;
    ram_cell[     498] = 32'hb15b0d5d;
    ram_cell[     499] = 32'h8897b0be;
    ram_cell[     500] = 32'hf928899c;
    ram_cell[     501] = 32'h99c19790;
    ram_cell[     502] = 32'hba6d862d;
    ram_cell[     503] = 32'h7ea51af4;
    ram_cell[     504] = 32'he752a496;
    ram_cell[     505] = 32'h08a710c7;
    ram_cell[     506] = 32'hc4dcc5a4;
    ram_cell[     507] = 32'hafa121ba;
    ram_cell[     508] = 32'h34fab601;
    ram_cell[     509] = 32'hcc0788b1;
    ram_cell[     510] = 32'h5a72f259;
    ram_cell[     511] = 32'h9dc8d3da;
    // src matrix B
    ram_cell[     512] = 32'h45fbb093;
    ram_cell[     513] = 32'hc863e305;
    ram_cell[     514] = 32'had04c01b;
    ram_cell[     515] = 32'hdd079c15;
    ram_cell[     516] = 32'h6bbf6513;
    ram_cell[     517] = 32'h66d47461;
    ram_cell[     518] = 32'h0dd6ff8e;
    ram_cell[     519] = 32'he9cab205;
    ram_cell[     520] = 32'hef611668;
    ram_cell[     521] = 32'hf4061912;
    ram_cell[     522] = 32'hbaa4a638;
    ram_cell[     523] = 32'h5f852dfa;
    ram_cell[     524] = 32'heeebfc25;
    ram_cell[     525] = 32'h04ce8a7c;
    ram_cell[     526] = 32'h09a3438e;
    ram_cell[     527] = 32'h532584c2;
    ram_cell[     528] = 32'hdb48cef5;
    ram_cell[     529] = 32'h48bc370b;
    ram_cell[     530] = 32'hee994a50;
    ram_cell[     531] = 32'hc1def925;
    ram_cell[     532] = 32'h1d7e8d48;
    ram_cell[     533] = 32'h2e770fab;
    ram_cell[     534] = 32'hac1e968b;
    ram_cell[     535] = 32'hd1ae8e2d;
    ram_cell[     536] = 32'hca1f0afa;
    ram_cell[     537] = 32'he41c3203;
    ram_cell[     538] = 32'ha1ba83b8;
    ram_cell[     539] = 32'h497efccc;
    ram_cell[     540] = 32'h6ee7b15e;
    ram_cell[     541] = 32'h851a3948;
    ram_cell[     542] = 32'h962bae50;
    ram_cell[     543] = 32'h0f0565cf;
    ram_cell[     544] = 32'h7b79e63d;
    ram_cell[     545] = 32'he1ec6b82;
    ram_cell[     546] = 32'h1483d926;
    ram_cell[     547] = 32'hece9b65c;
    ram_cell[     548] = 32'h10804931;
    ram_cell[     549] = 32'he9781068;
    ram_cell[     550] = 32'h7df4a173;
    ram_cell[     551] = 32'h145e8f00;
    ram_cell[     552] = 32'h0d7ccc6b;
    ram_cell[     553] = 32'he16eb293;
    ram_cell[     554] = 32'h7b2b0547;
    ram_cell[     555] = 32'he1b69fbd;
    ram_cell[     556] = 32'h53e6e51e;
    ram_cell[     557] = 32'h10d9dd06;
    ram_cell[     558] = 32'ha29d53fb;
    ram_cell[     559] = 32'h7fe631e7;
    ram_cell[     560] = 32'h9b4f087c;
    ram_cell[     561] = 32'hbe49af86;
    ram_cell[     562] = 32'h7f4c7cd6;
    ram_cell[     563] = 32'hd9af53f5;
    ram_cell[     564] = 32'hb7f6e0f5;
    ram_cell[     565] = 32'h6a065ef8;
    ram_cell[     566] = 32'h150ac737;
    ram_cell[     567] = 32'h1aae53dd;
    ram_cell[     568] = 32'hf4f0f094;
    ram_cell[     569] = 32'hbdf07d1b;
    ram_cell[     570] = 32'h74a298e6;
    ram_cell[     571] = 32'he1bd09af;
    ram_cell[     572] = 32'haf803bad;
    ram_cell[     573] = 32'h23981365;
    ram_cell[     574] = 32'hbcab1e46;
    ram_cell[     575] = 32'h127b8b03;
    ram_cell[     576] = 32'h60551211;
    ram_cell[     577] = 32'h838cfe5a;
    ram_cell[     578] = 32'h2bcb3aeb;
    ram_cell[     579] = 32'h411d866b;
    ram_cell[     580] = 32'h82858ba2;
    ram_cell[     581] = 32'h26fe3b4b;
    ram_cell[     582] = 32'hfa6f475e;
    ram_cell[     583] = 32'h0163bd1e;
    ram_cell[     584] = 32'h6d7e8ef7;
    ram_cell[     585] = 32'h697a832c;
    ram_cell[     586] = 32'h99539099;
    ram_cell[     587] = 32'h884382a5;
    ram_cell[     588] = 32'h8881e004;
    ram_cell[     589] = 32'h636b0023;
    ram_cell[     590] = 32'h6b32fd4e;
    ram_cell[     591] = 32'h1847b6ef;
    ram_cell[     592] = 32'h0ee8f22b;
    ram_cell[     593] = 32'h1b7eefc4;
    ram_cell[     594] = 32'hdab9a869;
    ram_cell[     595] = 32'h51266e59;
    ram_cell[     596] = 32'h6e5e8ba2;
    ram_cell[     597] = 32'hbb320387;
    ram_cell[     598] = 32'h0e272af9;
    ram_cell[     599] = 32'hcc290d56;
    ram_cell[     600] = 32'h299bb30d;
    ram_cell[     601] = 32'h3d741712;
    ram_cell[     602] = 32'h4c240790;
    ram_cell[     603] = 32'hd12fe580;
    ram_cell[     604] = 32'h5773f73c;
    ram_cell[     605] = 32'h1b30ae77;
    ram_cell[     606] = 32'h62153a9b;
    ram_cell[     607] = 32'h4dd2c52d;
    ram_cell[     608] = 32'h3b9a79a8;
    ram_cell[     609] = 32'h22e6c0fb;
    ram_cell[     610] = 32'h302aad5f;
    ram_cell[     611] = 32'hb4323bec;
    ram_cell[     612] = 32'h8ef37e7c;
    ram_cell[     613] = 32'h0b28a1b5;
    ram_cell[     614] = 32'hd25be998;
    ram_cell[     615] = 32'h9ab850c5;
    ram_cell[     616] = 32'h4f07579d;
    ram_cell[     617] = 32'h63f8697c;
    ram_cell[     618] = 32'hb416b9b0;
    ram_cell[     619] = 32'h4917046f;
    ram_cell[     620] = 32'h071eef5f;
    ram_cell[     621] = 32'h3e6689f1;
    ram_cell[     622] = 32'h05372976;
    ram_cell[     623] = 32'h0cf322bb;
    ram_cell[     624] = 32'h95907d50;
    ram_cell[     625] = 32'h72476793;
    ram_cell[     626] = 32'h320b9d4a;
    ram_cell[     627] = 32'h975a7cf6;
    ram_cell[     628] = 32'h1579f846;
    ram_cell[     629] = 32'h6bf250bb;
    ram_cell[     630] = 32'heeae01d5;
    ram_cell[     631] = 32'h25a15c66;
    ram_cell[     632] = 32'h839683a1;
    ram_cell[     633] = 32'h2d029132;
    ram_cell[     634] = 32'h5a2c2281;
    ram_cell[     635] = 32'h2c887b00;
    ram_cell[     636] = 32'hc94533f6;
    ram_cell[     637] = 32'h78508abe;
    ram_cell[     638] = 32'h5fe5ae86;
    ram_cell[     639] = 32'he580814e;
    ram_cell[     640] = 32'hcd06d6db;
    ram_cell[     641] = 32'h912676ea;
    ram_cell[     642] = 32'h9f3b363d;
    ram_cell[     643] = 32'h0e96376e;
    ram_cell[     644] = 32'ha147b195;
    ram_cell[     645] = 32'h12a98a5d;
    ram_cell[     646] = 32'h508ecb19;
    ram_cell[     647] = 32'hbd729370;
    ram_cell[     648] = 32'h39a6c099;
    ram_cell[     649] = 32'h7ed64243;
    ram_cell[     650] = 32'h1135d57f;
    ram_cell[     651] = 32'h7562d9e0;
    ram_cell[     652] = 32'h48bc433d;
    ram_cell[     653] = 32'hcd7e224d;
    ram_cell[     654] = 32'h926fbac5;
    ram_cell[     655] = 32'h282a7faa;
    ram_cell[     656] = 32'h8d2af208;
    ram_cell[     657] = 32'h441ff440;
    ram_cell[     658] = 32'hcf7efd4b;
    ram_cell[     659] = 32'h2670bcd0;
    ram_cell[     660] = 32'h8b9e0d51;
    ram_cell[     661] = 32'ha085c219;
    ram_cell[     662] = 32'h073a4870;
    ram_cell[     663] = 32'he50b705c;
    ram_cell[     664] = 32'haa540e28;
    ram_cell[     665] = 32'h243d956c;
    ram_cell[     666] = 32'hb0bd9d28;
    ram_cell[     667] = 32'h9710a762;
    ram_cell[     668] = 32'ha27accb1;
    ram_cell[     669] = 32'he060b2d0;
    ram_cell[     670] = 32'hf88d6f6d;
    ram_cell[     671] = 32'had29b4dc;
    ram_cell[     672] = 32'hfb0ede70;
    ram_cell[     673] = 32'hdf7f1512;
    ram_cell[     674] = 32'h0178cafc;
    ram_cell[     675] = 32'h6b46b61b;
    ram_cell[     676] = 32'h6da7d4c7;
    ram_cell[     677] = 32'hf5d47d24;
    ram_cell[     678] = 32'h9408a139;
    ram_cell[     679] = 32'he91a2912;
    ram_cell[     680] = 32'h7232b853;
    ram_cell[     681] = 32'hb25be49d;
    ram_cell[     682] = 32'hb162f411;
    ram_cell[     683] = 32'h499b8fc4;
    ram_cell[     684] = 32'hd25b3f71;
    ram_cell[     685] = 32'h6870c704;
    ram_cell[     686] = 32'he1b55027;
    ram_cell[     687] = 32'h983c164b;
    ram_cell[     688] = 32'h5c597840;
    ram_cell[     689] = 32'h0f85a26a;
    ram_cell[     690] = 32'h30164325;
    ram_cell[     691] = 32'h0809a682;
    ram_cell[     692] = 32'hc3d7919e;
    ram_cell[     693] = 32'h9ebae8a0;
    ram_cell[     694] = 32'h75c590d2;
    ram_cell[     695] = 32'h5263c656;
    ram_cell[     696] = 32'h65525d38;
    ram_cell[     697] = 32'h5483b3bd;
    ram_cell[     698] = 32'heff53260;
    ram_cell[     699] = 32'he892829a;
    ram_cell[     700] = 32'hd632f2c5;
    ram_cell[     701] = 32'hc30a167f;
    ram_cell[     702] = 32'h24315d0d;
    ram_cell[     703] = 32'ha8b931f4;
    ram_cell[     704] = 32'h88a90edc;
    ram_cell[     705] = 32'h7fc7fa48;
    ram_cell[     706] = 32'h432482ca;
    ram_cell[     707] = 32'h47c1b174;
    ram_cell[     708] = 32'h4c1c0388;
    ram_cell[     709] = 32'hda7e9fce;
    ram_cell[     710] = 32'h78fddc99;
    ram_cell[     711] = 32'hb853bf5b;
    ram_cell[     712] = 32'h094debfe;
    ram_cell[     713] = 32'hbfddc135;
    ram_cell[     714] = 32'h8d279b5b;
    ram_cell[     715] = 32'h89b8c0a4;
    ram_cell[     716] = 32'h45745085;
    ram_cell[     717] = 32'h0d5c43cb;
    ram_cell[     718] = 32'hd43ad07e;
    ram_cell[     719] = 32'he996e3dd;
    ram_cell[     720] = 32'hf8cda506;
    ram_cell[     721] = 32'h46e7996b;
    ram_cell[     722] = 32'h6cd77c60;
    ram_cell[     723] = 32'h345835f3;
    ram_cell[     724] = 32'he18b8f3b;
    ram_cell[     725] = 32'h9f14387b;
    ram_cell[     726] = 32'h7d9e0e34;
    ram_cell[     727] = 32'hebca4553;
    ram_cell[     728] = 32'h3ffee786;
    ram_cell[     729] = 32'h23b9c390;
    ram_cell[     730] = 32'hd18e07e9;
    ram_cell[     731] = 32'hbba0f62e;
    ram_cell[     732] = 32'h995c1b35;
    ram_cell[     733] = 32'hee0ee420;
    ram_cell[     734] = 32'h16e481b5;
    ram_cell[     735] = 32'h54dc52d3;
    ram_cell[     736] = 32'h8188dd5c;
    ram_cell[     737] = 32'he12d53b2;
    ram_cell[     738] = 32'hd2c9b837;
    ram_cell[     739] = 32'h0c513105;
    ram_cell[     740] = 32'h79611cab;
    ram_cell[     741] = 32'h88bb79c9;
    ram_cell[     742] = 32'h41043728;
    ram_cell[     743] = 32'h474d17b4;
    ram_cell[     744] = 32'h0e313366;
    ram_cell[     745] = 32'h6a836011;
    ram_cell[     746] = 32'ha9361388;
    ram_cell[     747] = 32'h8932e69f;
    ram_cell[     748] = 32'hba29c360;
    ram_cell[     749] = 32'h91e9a2de;
    ram_cell[     750] = 32'h7b835b35;
    ram_cell[     751] = 32'hfbcae232;
    ram_cell[     752] = 32'h24a0f2f5;
    ram_cell[     753] = 32'h8e2d3455;
    ram_cell[     754] = 32'h85e3ff51;
    ram_cell[     755] = 32'h0b4e71a7;
    ram_cell[     756] = 32'hd66141f0;
    ram_cell[     757] = 32'h14fdec60;
    ram_cell[     758] = 32'h6aa79824;
    ram_cell[     759] = 32'h1e628f44;
    ram_cell[     760] = 32'h0b8ea51b;
    ram_cell[     761] = 32'h79f695db;
    ram_cell[     762] = 32'h44e0211d;
    ram_cell[     763] = 32'hb243982d;
    ram_cell[     764] = 32'h823c0907;
    ram_cell[     765] = 32'h59c969cb;
    ram_cell[     766] = 32'h65c5a0a6;
    ram_cell[     767] = 32'hb31d1bc2;
end

endmodule

